module lab2 (
	CLOCK_50,

	HEX0,							
	HEX1,								
	HEX2,
	HEX3,
	HEX4,
	HEX5,

	KEY,

	LEDR,

	SW,

	HPS_DDR3_ADDR,
	HPS_DDR3_BA,
	HPS_DDR3_CAS_N,
	HPS_DDR3_CKE,
	HPS_DDR3_CK_N,
	HPS_DDR3_CK_P,
	HPS_DDR3_CS_N,
	HPS_DDR3_RESET_N,
	HPS_DDR3_RZQ,
	HPS_DDR3_WE_N, 
	
	HPS_DDR3_DM,
	HPS_DDR3_DQ,
	HPS_DDR3_DQS_N,
	HPS_DDR3_DQS_P,
	HPS_DDR3_ODT,
	HPS_DDR3_RAS_N,
	
	
	DRAM_CLK
);

	input CLOCK_50;
	output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
	input [3:0] KEY;
	output [9:0] LEDR;
	input [9:0] SW;

	output [14:0] HPS_DDR3_ADDR;
	output [2:0] HPS_DDR3_BA;
	output HPS_DDR3_CAS_N;
	output HPS_DDR3_CKE;
	output HPS_DDR3_CK_N;
	output HPS_DDR3_CK_P;
	output HPS_DDR3_CS_N;
	output [3:0] HPS_DDR3_DM;
	inout [31:0] HPS_DDR3_DQ;
	inout [3:0] HPS_DDR3_DQS_N;
	inout [3:0] HPS_DDR3_DQS_P;
	output HPS_DDR3_ODT;
	output HPS_DDR3_RAS_N;
	output HPS_DDR3_RESET_N;
	input HPS_DDR3_RZQ;
	output HPS_DDR3_WE_N;
	
	input DRAM_CLK;
	wire [31:0] INT_IN;
	//assign INT_IN= 255;
	wire [31:0] hex3_hex0;
	wire [15:0] hex5_hex4;
	wire [9:0] ledR;

//	assign HEX0 = ~hex3_hex0[6:0];
//	assign HEX1 = ~hex3_hex0[14:8];
//	assign HEX2 = ~hex3_hex0[22:16];
//	assign HEX3 = ~hex3_hex0[30:24];
//	assign HEX4 = ~hex5_hex4[6:0];
//	assign HEX5 = ~hex5_hex4[14:8];
	
	assign LEDR = {2'b0, INT_IN[31:24]}; 
	
	display_hex h0(INT_IN[3:0], HEX0);
	display_hex h1(INT_IN[7:4], HEX1);
	display_hex h2(INT_IN[11:8], HEX2);
	display_hex h3(INT_IN[15:12], HEX3);
	display_hex h4(INT_IN[19:16], HEX4);
	display_hex h5(INT_IN[23:20], HEX5);

    mysystem u0 (
        //.hex3_0bus_export       (hex3_hex0),       //        hex3_0bus.export
        //.hex5_4bus_export       (hex5_hex4),       //        hex5_4bus.export
        .memory_mem_a           (HPS_DDR3_ADDR),           //           memory.mem_a
        .memory_mem_ba          (HPS_DDR3_BA),          //                 .mem_ba
        .memory_mem_ck          (HPS_DDR3_CK_P),          //                 .mem_ck
        .memory_mem_ck_n        (HPS_DDR3_CK_N),        //                 .mem_ck_n
        .memory_mem_cke         (HPS_DDR3_CKE),         //                 .mem_cke
        .memory_mem_cs_n        (HPS_DDR3_CS_N),        //                 .mem_cs_n
        .memory_mem_ras_n       (HPS_DDR3_RAS_N),       //                 .mem_ras_n
        .memory_mem_cas_n       (HPS_DDR3_CAS_N),       //                 .mem_cas_n
        .memory_mem_we_n        (HPS_DDR3_WE_N),        //                 .mem_we_n
        .memory_mem_reset_n     (HPS_DDR3_RESET_N),     //                 .mem_reset_n
        .memory_mem_dq          (HPS_DDR3_DQ),          //                 .mem_dq
        .memory_mem_dqs         (HPS_DDR3_DQS_P),         //                 .mem_dqs
        .memory_mem_dqs_n       (HPS_DDR3_DQS_N),       //                 .mem_dqs_n
        .memory_mem_odt         (HPS_DDR3_ODT),         //                 .mem_odt
        .memory_mem_dm          (HPS_DDR3_DM),          //                 .mem_dm
        .memory_oct_rzqin       (HPS_DDR3_RZQ),       //                 .oct_rzqin
        .pushbutton_export      ({~KEY[3:1], 1'b0}),      //       pushbutton.export
        .sdram_clk_clk          (DRAM_CLK),          //        sdram_clk.clk
        .system_ref_clk_clk     (CLOCK_50),     //   system_ref_clk.clk
        .system_ref_reset_reset (~KEY[0]), // system_ref_reset.reset
        .to_hex_to_led_readdata (INT_IN)  //    to_hex_to_led.readdata
    );


endmodule